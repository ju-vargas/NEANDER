library verilog;
use verilog.vl_types.all;
entity decod_vlg_check_tst is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        d3              : in     vl_logic;
        d4              : in     vl_logic;
        d5              : in     vl_logic;
        d6              : in     vl_logic;
        d7              : in     vl_logic;
        d8              : in     vl_logic;
        d9              : in     vl_logic;
        d10             : in     vl_logic;
        d11             : in     vl_logic;
        d12             : in     vl_logic;
        d13             : in     vl_logic;
        d14             : in     vl_logic;
        d15             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end decod_vlg_check_tst;
