library verilog;
use verilog.vl_types.all;
entity neander_top_vlg_vec_tst is
end neander_top_vlg_vec_tst;
