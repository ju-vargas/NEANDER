library verilog;
use verilog.vl_types.all;
entity name_top_vlg_vec_tst is
end name_top_vlg_vec_tst;
