library verilog;
use verilog.vl_types.all;
entity NeanderMain_vlg_vec_tst is
end NeanderMain_vlg_vec_tst;
