library verilog;
use verilog.vl_types.all;
entity ula16_vlg_vec_tst is
end ula16_vlg_vec_tst;
