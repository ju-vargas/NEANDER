library verilog;
use verilog.vl_types.all;
entity uctop_vlg_vec_tst is
end uctop_vlg_vec_tst;
